module hello_module;
    initial begin
        $display("Hello");
    end
endmodule
