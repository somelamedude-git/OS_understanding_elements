module not_gate(input wire a, output wire y);
    not(y, a);
endmodule
