module not_gate(input reg a, output wire y);
    not(y, a);
endmodule
