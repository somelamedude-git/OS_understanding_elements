module or_gate(input wire a, input wire b, output wire y);
    or(y,a,b);
endmodule
