module and_gate(input wire a, input wire b, output wire y);
    and(y,a,b);
endmodule
